// module memory_controller.v

// WORK_STATE: 

// load datas [head_addr, head_addr + length) from memory

