// module instruction_fetcher.v

// use module_Decoder to decode the instruction
// interact with Branch_Predictor to get the next PC
// interact with ICache to get the instruction at PC
// interact with Dispatcher to send the instruction to Dispatcher
// FLUSH: when predict goes wrong




