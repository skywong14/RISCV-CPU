// module CDB.v